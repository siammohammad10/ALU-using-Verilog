// =========================== TESTBENCH: AND =========================== //
`timescale 1ns / 1ps
`include "and.v"

module tb_and;
    reg [7:0] opA, opB;
    wire [7:0] result;

    AND uut(
        .result(result),
        .opA(opA), .opB(opB)
    );

    initial begin
        $display("Testing AND");

        // Example test case
        opA = 8'd15;
        opB = 8'd3;
        #1 $display("opA = %d, opB = %d, result = %d", opA, opB, result);
        
        // Additional test cases can be added here
        $finish;
    end
endmodule

// iverilog -o tb_and.vvp tb_and.v
// vvp tb_and.vvp

