// =========================== TESTBENCH: XOR =========================== //
`timescale 1ns / 1ps
`include "xor.v"

module tb_xor;
    reg [7:0] opA, opB;
    wire [7:0] result;

    XOR uut(
        .result(result),
        .opA(opA), .opB(opB)
    );

    initial begin
        $display("Testing XOR");

        // Example test case
        opA = 8'd15;
        opB = 8'd3;
        #1 $display("opA = %d, opB = %d, result = %d", opA, opB, result);
        
        // Additional test cases can be added here
        $finish;
    end
endmodule

// iverilog -o tb_xor.vvp tb_xor.v
// vvp tb_xor.vvp
