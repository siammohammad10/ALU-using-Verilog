// =========================== TESTBENCH: SHIFT_RIGHT =========================== //

`timescale 1ns / 1ps
`include "shift_right.v"

module tb_shift_right;
    reg [7:0] op;
    wire [7:0] result;

    SHIFT_RIGHT uut(
        .result(result),
        .op(op)
    );

    initial begin
        $display("Testing SHIFT_RIGHT");

        // Example test case
        op = 8'd15; // 00001111
        #10 $display("op = %b, result = %b", op, result); // Expected: 00000111

        op = 8'b00000001;
        #10 $display("op = %b, result = %b", op, result); // Expected: 00000000

        $finish;
    end
endmodule

// iverilog -o tb_shift_right.vvp tb_shift_right.v
// vvp tb_shift_right.vvp
